`timescale 1ns / 1ps 
`define TASK1_HANDLER_ENT 32'h800010e8
`define TASK1_DELETE 32'h80001310

`define IRQ_HANDLE_ENT 32'h80007400
`define PROCESSED_SRC_END 32'h800075e4 // -4

`define SEMAPHORE_TAKE_ENT 32'h8000338c
`define SEMAPHORE_TAKE_RET 32'h800034b8 // -4
`define SEMAPHORE_GIVE_ENT 32'h80002cc4
`define SEMAPHORE_GIVE_RET 32'h80002d74 // -4

`define ENTER_CRITICAL_ENT 32'h80004dc0
`define ENTER_CRITICAL_RET 32'h80004de8
`define EXIT_CRITICAL_ENT 32'h80004dec
`define EXIT_CRITICAL_RET 32'h80004e28

/*
`define IRQ_HANDLE_END 32'h8000748c
`define HANDLE_ASYNC_ENT 32'h8000749c
`define HANDLE_ASYNC_END 32'h80007504
`define TASK_INCR_ENT 32'h80004410
`define TASK_INCR_RET 32'h80004124 // part.0 return (part.0 => scheduler is not suspended)
`define CONTXT_SW_ENT 32'h8000444c
`define CONTXT_SW_RET 32'h8000451c
`define PROCESSED_SRC_ENT 32'h80007558
*/
